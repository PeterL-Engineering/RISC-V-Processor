module datapath(
    input logic clk,
    input logic reset,
    input logic 
)

endmodule